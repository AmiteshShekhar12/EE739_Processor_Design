library ieee;
use ieee.std_logic_1164.all;

entity In_Order_2_Way is
end entity;