library ieee;
use ieee.std_logic_1164.all;

entity MUX_2_3bit  is
  port (IN_0, IN_1: in std_logic_vector(2 downto 0);
			S : in std_logic;
			Y: out std_logic_vector(2 downto 0));
end entity MUX_2_3bit;

architecture Struct of MUX_2_3bit is
begin
bit_3_1 : for i in 0 to 2 generate 
		Y(i) <= (IN_0(i) AND (NOT S)) OR (IN_1(i) AND S);
end generate ;
end Struct;