--library ieee;
--use ieee.std_logic_1164.all;
--
--entity serial_shift_reg_rs is
--	port (